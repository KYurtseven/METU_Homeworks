`timescale 1ns / 1ps
module ALU(
input [3:0] A, 
input [3:0] B, 
input [3:0] ALUop, 
output reg [3:0] C, 
output reg [3:0] Cond // Z,N,C,V
    );
//
//Write your code below
//
	
endmodule