    CONSTANT MaxMem   : NATURAL := 16#FF#;  
    TYPE     MemArrayT IS ARRAY(0 TO MaxMem-1) OF ByteT;
    VARIABLE Mem  : MemArrayT
            :=  (-- program
                 3=>"01100000",  2=>"00000000",  1=>"00000000",  0=>"00000000",
                 7=>"01000100",  6=>"00100000",  5=>"00000000",  4=>"00110010",
                11=>"10000110", 10=>"10000001",  9=>"00000000",  8=>"00000000",
                15=>"10000110", 14=>"10100001", 13=>"00000000", 12=>"00000100",
                19=>"01000100", 18=>"01000000", 17=>"00000000", 16=>"00111111",
                23=>"10001000", 22=>"01000001", 21=>"00000000", 20=>"00000000",
              -- data
                51=>"00110011", 50=>"00001111", 49=>"11110000", 48=>"11001100",
                55=>"00110011", 54=>"00001111", 53=>"11110000", 52=>"11001100",
                OTHERS => "00000000");

